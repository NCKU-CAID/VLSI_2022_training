`include "DRAM.sv"

module DRAM_wrapper (
);

	

endmodule
